module zero_detection(
	input [31:0] result,
	output zero_bit
);
	nor nor0(zero_bit,
		result[31],
		result[30],
		result[29],
		result[28],
		result[27],
		result[26],
		result[25],
		result[24],
		result[23],
		result[22],
		result[21],
		result[20],
		result[19],
		result[18],
		result[17],
		result[16],
		result[15],
		result[14],
		result[13],
		result[12],
		result[11],
		result[10],
		result[9],
		result[8],
		result[7],
		result[6],
		result[5],
		result[4],
		result[3],
		result[2],
		result[1],
		result[0]);

endmodule
